module ROM (
    input wire edit,          // 编程模式信号
    input wire [7:0] unit,    // 代码位置
    input wire [7:0] code,    // 代码
    input wire send,          // 发送程序信号
    input wire clk,           // 时钟信号
    input wire rst,           // 复位信号
    input wire [7:0] address, // 地址输入
    output reg [31:0] opcode  // 当前输出的机器码
);

localparam IMM1 = 8'b10000000;
localparam IMM2 = 8'b01000000;
localparam MOV  = 8'b01000000;
localparam JMP  = 8'b10000000;
localparam PUSH = 8'b01000000;
localparam POP  = 8'b01000000;
localparam TO   = 8'b00000000;
localparam ADD = 8'b00000000;
localparam SUB = 8'b00000001;
localparam AND = 8'b00000010;
localparam OR  = 8'b00000011;
localparam NOT = 8'b00000100;
localparam XOR = 8'b00000101;
localparam SHL = 8'b00000110;
localparam SHR = 8'b00000111;
localparam MUL = 8'b00001000;
localparam DIV = 8'b00001001;
localparam MOD = 8'b00001010;
localparam NULL    = 8'b00000000;
localparam REG0    = 8'b00000000;
localparam REG1    = 8'b00000001;
localparam REG2    = 8'b00000010;
localparam REG3    = 8'b00000011;
localparam REG4    = 8'b00000100;
localparam REG5    = 8'b00000101;
localparam RAM     = 8'b00010000;
localparam REG_RAM = 8'b00010001;
localparam STACK   = 8'b00010010;
localparam COUNTER = 8'b00000110;
localparam INPUT   = 8'b00000111;
localparam OUTPUT  = 8'b00000111;
localparam IF_EQUAL            = 8'b10000000;
localparam IF_NOT_EQUAL        = 8'b10000001;
localparam IF_LESS             = 8'b10000010;
localparam IF_LESS_OR_EQUAL    = 8'b10000011;
localparam IF_GREATER          = 8'b10010000;
localparam IF_GREATER_OR_EQUAL = 8'b10010001;
localparam CALL = 8'b00110000;
localparam RET  = 8'b00110001;
localparam HALT = 8'b00110010;

reg [7:0] memory [0:255];     // 16*16 = 256个8位机器码

/**
CONST IO_NUM 32
IMM1|MOV         0           TO          REG_RAM    # REG_RAM置0
# 循环INPUT:
LABEL CIRCLE_I
IMM2|IF_EQUAL    REG_RAM     IO_NUM      DATA_O     # 如果REG_RAM=IO_NUM，跳转到DATA_O
MOV              INPUT       TO          RAM        # RAM <- INPUT
IMM2|ADD         REG_RAM     1           REG_RAM    # REG_RAM++
IMM2|JMP         TO          CIRCLE_I    COUNTER    # 跳转到CIRCLE_I
# 循环OUTPUT:
LABEL DATA_O
IMM1|MOV         0           TO          REG_RAM    # REG_RAM置0
LABEL CIRCLE_O
IMM2|IF_EQUAL    REG_RAM     IO_NUM      END        # 如果REG_RAM=IO_NUM，跳转到END结束
MOV              RAM         TO          OUTPUT     # OUTPUT <- RAM
IMM2|ADD         REG_RAM     1           REG_RAM    # REG_RAM++
IMM1|MOV         CIRCLE_O    TO          COUNTER    # COUNTER <- CIRCLE_O
LABEL END
**/
localparam IO_NUM = 8'b00100000; // 每次读32个
always @(posedge clk or posedge rst) begin
    if (rst) begin // 这是ROM (BIOS)
        memory[0]  <= (IMM1 | MOV);               // 0: IMM1 | MOV
        memory[1]  <= 8'b00000000;              // 1: 0
        memory[2]  <= TO;                       // 2: TO
        memory[3]  <= REG_RAM;                  // 3: REG_RAM
        // 循环INPUT
        memory[4]  <= IMM2 | IF_EQUAL;          // 4: IMM2 | IF_EQUAL
        memory[5]  <= REG_RAM;                  // 5: REG_RAM
        memory[6]  <= IO_NUM;                   // 6: IO_NUM
        memory[7]  <= 8'b00010100;              // 7: DATA_O: 20
        memory[8]  <= MOV;                      // 8: MOV
        memory[9]  <= INPUT;                    // 9: INPUT
        memory[10] <= TO;                       // 10: TO
        memory[11] <= RAM;                      // 11: RAM
        memory[12] <= IMM2 | ADD;               // 12: IMM2 | ADD
        memory[13] <= REG_RAM;                  // 13: REG_RAM
        memory[14] <= 8'b00000001;              // 14: 1
        memory[15] <= REG_RAM;                  // 15: REG_RAM
        memory[16] <= IMM2 | JMP;               // 16: IMM2 | JMP
        memory[17] <= TO;                       // 17: TO
        memory[18] <= 8'b00000100;              // 18: CIRCLE_I: 4
        memory[19] <= COUNTER;                  // 19: COUNTER
        // 循环OUTPUT
        memory[20] <= IMM1 | MOV;               // 20: IMM1 | MOV
        memory[21] <= 8'b00000000;              // 21: 0
        memory[22] <= TO;                       // 22: TO
        memory[23] <= REG_RAM;                  // 23: REG_RAM
        memory[24] <= IMM2 | IF_EQUAL;          // 24: IMM2 | IF_EQUAL
        memory[25] <= REG_RAM;                  // 25: REG_RAM
        memory[26] <= IO_NUM;                   // 26: IO_NUM
        memory[27] <= 8'b00101000;              // 27: END: 40
        memory[28] <= MOV;                      // 28: MOV
        memory[29] <= RAM;                      // 29: RAM
        memory[30] <= TO;                       // 30: TO
        memory[31] <= OUTPUT;                   // 31: OUTPUT
        memory[32] <= IMM2 | ADD;               // 32: IMM2 | ADD
        memory[33] <= REG_RAM;                  // 33: REG_RAM
        memory[34] <= 8'b00000001;              // 34: 1
        memory[35] <= REG_RAM;                  // 35: REG_RAM
        memory[36] <= IMM1 | MOV;               // 36: IMM1 | MOV
        memory[37] <= 8'b00000100;              // 37: CIRCLE_O: 4
        memory[38] <= TO;                       // 38: TO
        memory[39] <= COUNTER;                  // 39: COUNTER
        memory[40] <= HALT;                     // 40: HALT
        memory[41] <= 8'b00000000;
        memory[42] <= 8'b00000000;
        memory[43] <= 8'b00000000;
        memory[44] <= 8'b00000000;
        memory[45] <= 8'b00000000;
        memory[46] <= 8'b00000000;
        memory[47] <= 8'b00000000;
        memory[48] <= 8'b00000000;
        memory[49] <= 8'b00000000;
        memory[50] <= 8'b00000000;
        memory[51] <= 8'b00000000;
        memory[52] <= 8'b00000000;
        memory[53] <= 8'b00000000;
        memory[54] <= 8'b00000000;
        memory[55] <= 8'b00000000;
        memory[56] <= 8'b00000000;
        memory[57] <= 8'b00000000;
        memory[58] <= 8'b00000000;
        memory[59] <= 8'b00000000;
        memory[60] <= 8'b00000000;
        memory[61] <= 8'b00000000;
        memory[62] <= 8'b00000000;
        memory[63] <= 8'b00000000;
        memory[64] <= 8'b00000000;
        memory[65] <= 8'b00000000;
        memory[66] <= 8'b00000000;
        memory[67] <= 8'b00000000;
        memory[68] <= 8'b00000000;
        memory[69] <= 8'b00000000;
        memory[70] <= 8'b00000000;
        memory[71] <= 8'b00000000;
        memory[72] <= 8'b00000000;
        memory[73] <= 8'b00000000;
        memory[74] <= 8'b00000000;
        memory[75] <= 8'b00000000;
        memory[76] <= 8'b00000000;
        memory[77] <= 8'b00000000;
        memory[78] <= 8'b00000000;
        memory[79] <= 8'b00000000;
        memory[80] <= 8'b00000000;
        memory[81] <= 8'b00000000;
        memory[82] <= 8'b00000000;
        memory[83] <= 8'b00000000;
        memory[84] <= 8'b00000000;
        memory[85] <= 8'b00000000;
        memory[86] <= 8'b00000000;
        memory[87] <= 8'b00000000;
        memory[88] <= 8'b00000000;
        memory[89] <= 8'b00000000;
        memory[90] <= 8'b00000000;
        memory[91] <= 8'b00000000;
        memory[92] <= 8'b00000000;
        memory[93] <= 8'b00000000;
        memory[94] <= 8'b00000000;
        memory[95] <= 8'b00000000;
        memory[96] <= 8'b00000000;
        memory[97] <= 8'b00000000;
        memory[98] <= 8'b00000000;
        memory[99] <= 8'b00000000;
        memory[100] <= 8'b00000000;
        memory[101] <= 8'b00000000;
        memory[102] <= 8'b00000000;
        memory[103] <= 8'b00000000;
        memory[104] <= 8'b00000000;
        memory[105] <= 8'b00000000;
        memory[106] <= 8'b00000000;
        memory[107] <= 8'b00000000;
        memory[108] <= 8'b00000000;
        memory[109] <= 8'b00000000;
        memory[110] <= 8'b00000000;
        memory[111] <= 8'b00000000;
        memory[112] <= 8'b00000000;
        memory[113] <= 8'b00000000;
        memory[114] <= 8'b00000000;
        memory[115] <= 8'b00000000;
        memory[116] <= 8'b00000000;
        memory[117] <= 8'b00000000;
        memory[118] <= 8'b00000000;
        memory[119] <= 8'b00000000;
        memory[120] <= 8'b00000000;
        memory[121] <= 8'b00000000;
        memory[122] <= 8'b00000000;
        memory[123] <= 8'b00000000;
        memory[124] <= 8'b00000000;
        memory[125] <= 8'b00000000;
        memory[126] <= 8'b00000000;
        memory[127] <= 8'b00000000;
        memory[128] <= 8'b00000000;
        memory[129] <= 8'b00000000;
        memory[130] <= 8'b00000000;
        memory[131] <= 8'b00000000;
        memory[132] <= 8'b00000000;
        memory[133] <= 8'b00000000;
        memory[134] <= 8'b00000000;
        memory[135] <= 8'b00000000;
        memory[136] <= 8'b00000000;
        memory[137] <= 8'b00000000;
        memory[138] <= 8'b00000000;
        memory[139] <= 8'b00000000;
        memory[140] <= 8'b00000000;
        memory[141] <= 8'b00000000;
        memory[142] <= 8'b00000000;
        memory[143] <= 8'b00000000;
        memory[144] <= 8'b00000000;
        memory[145] <= 8'b00000000;
        memory[146] <= 8'b00000000;
        memory[147] <= 8'b00000000;
        memory[148] <= 8'b00000000;
        memory[149] <= 8'b00000000;
        memory[150] <= 8'b00000000;
        memory[151] <= 8'b00000000;
        memory[152] <= 8'b00000000;
        memory[153] <= 8'b00000000;
        memory[154] <= 8'b00000000;
        memory[155] <= 8'b00000000;
        memory[156] <= 8'b00000000;
        memory[157] <= 8'b00000000;
        memory[158] <= 8'b00000000;
        memory[159] <= 8'b00000000;
        memory[160] <= 8'b00000000;
        memory[161] <= 8'b00000000;
        memory[162] <= 8'b00000000;
        memory[163] <= 8'b00000000;
        memory[164] <= 8'b00000000;
        memory[165] <= 8'b00000000;
        memory[166] <= 8'b00000000;
        memory[167] <= 8'b00000000;
        memory[168] <= 8'b00000000;
        memory[169] <= 8'b00000000;
        memory[170] <= 8'b00000000;
        memory[171] <= 8'b00000000;
        memory[172] <= 8'b00000000;
        memory[173] <= 8'b00000000;
        memory[174] <= 8'b00000000;
        memory[175] <= 8'b00000000;
        memory[176] <= 8'b00000000;
        memory[177] <= 8'b00000000;
        memory[178] <= 8'b00000000;
        memory[179] <= 8'b00000000;
        memory[180] <= 8'b00000000;
        memory[181] <= 8'b00000000;
        memory[182] <= 8'b00000000;
        memory[183] <= 8'b00000000;
        memory[184] <= 8'b00000000;
        memory[185] <= 8'b00000000;
        memory[186] <= 8'b00000000;
        memory[187] <= 8'b00000000;
        memory[188] <= 8'b00000000;
        memory[189] <= 8'b00000000;
        memory[190] <= 8'b00000000;
        memory[191] <= 8'b00000000;
        memory[192] <= 8'b00000000;
        memory[193] <= 8'b00000000;
        memory[194] <= 8'b00000000;
        memory[195] <= 8'b00000000;
        memory[196] <= 8'b00000000;
        memory[197] <= 8'b00000000;
        memory[198] <= 8'b00000000;
        memory[199] <= 8'b00000000;
        memory[200] <= 8'b00000000;
        memory[201] <= 8'b00000000;
        memory[202] <= 8'b00000000;
        memory[203] <= 8'b00000000;
        memory[204] <= 8'b00000000;
        memory[205] <= 8'b00000000;
        memory[206] <= 8'b00000000;
        memory[207] <= 8'b00000000;
        memory[208] <= 8'b00000000;
        memory[209] <= 8'b00000000;
        memory[210] <= 8'b00000000;
        memory[211] <= 8'b00000000;
        memory[212] <= 8'b00000000;
        memory[213] <= 8'b00000000;
        memory[214] <= 8'b00000000;
        memory[215] <= 8'b00000000;
        memory[216] <= 8'b00000000;
        memory[217] <= 8'b00000000;
        memory[218] <= 8'b00000000;
        memory[219] <= 8'b00000000;
        memory[220] <= 8'b00000000;
        memory[221] <= 8'b00000000;
        memory[222] <= 8'b00000000;
        memory[223] <= 8'b00000000;
        memory[224] <= 8'b00000000;
        memory[225] <= 8'b00000000;
        memory[226] <= 8'b00000000;
        memory[227] <= 8'b00000000;
        memory[228] <= 8'b00000000;
        memory[229] <= 8'b00000000;
        memory[230] <= 8'b00000000;
        memory[231] <= 8'b00000000;
        memory[232] <= 8'b00000000;
        memory[233] <= 8'b00000000;
        memory[234] <= 8'b00000000;
        memory[235] <= 8'b00000000;
        memory[236] <= 8'b00000000;
        memory[237] <= 8'b00000000;
        memory[238] <= 8'b00000000;
        memory[239] <= 8'b00000000;
        memory[240] <= 8'b00000000;
        memory[241] <= 8'b00000000;
        memory[242] <= 8'b00000000;
        memory[243] <= 8'b00000000;
        memory[244] <= 8'b00000000;
        memory[245] <= 8'b00000000;
        memory[246] <= 8'b00000000;
        memory[247] <= 8'b00000000;
        memory[248] <= 8'b00000000;
        memory[249] <= 8'b00000000;
        memory[250] <= 8'b00000000;
        memory[251] <= 8'b00000000;
        memory[252] <= 8'b00000000;
        memory[253] <= 8'b00000000;
        memory[254] <= 8'b00000000;
        memory[255] <= 8'b00000000;
        opcode <= 32'b0;
    end else if (edit & send)  begin
        memory[unit]  <= code;
    end else begin
        opcode <= {memory[address+3], memory[address+2], memory[address+1], memory[address]};
    end
end
endmodule
