module ROM (
    input wire clk,                     // 时钟信号
    input wire rst,                     // 复位信号
    input wire [7:0] address,           // 地址输入
    output reg [31:0] opcode,           // 当前输出的机器码

    input wire [7:0] monitor_inputs0,   // 监视寄存器输入0
    input wire [7:0] monitor_inputs1,   // 监视寄存器输入1
    input wire [7:0] monitor_inputs2,   // 监视寄存器输入2
    input wire [7:0] monitor_inputs3,   // 监视寄存器输入3
    input wire [7:0] monitor_inputs4,   // 监视寄存器输入4
    input wire [7:0] monitor_inputs5,   // 监视寄存器输入5
    input wire [7:0] monitor_inputs6,   // 监视寄存器输入6
    input wire [7:0] monitor_inputs7,   // 监视寄存器输入7
    input wire [7:0] monitor_inputs8,   // 监视寄存器输入8
    input wire [7:0] monitor_inputs9,   // 监视寄存器输入9
    input wire [7:0] monitor_inputs10,  // 监视寄存器输入10
    input wire [7:0] monitor_inputs11,  // 监视寄存器输入11
    input wire [7:0] monitor_inputs12,  // 监视寄存器输入12
    input wire [7:0] monitor_inputs13,  // 监视寄存器输入13
    input wire [7:0] monitor_inputs14,  // 监视寄存器输入14
    input wire [7:0] monitor_inputs15,  // 监视寄存器输入15
    output reg [7:0] monitor_outputs0,  // 监视输出0
    output reg [7:0] monitor_outputs1,  // 监视输出1
    output reg [7:0] monitor_outputs2,  // 监视输出2
    output reg [7:0] monitor_outputs3,  // 监视输出3
    output reg [7:0] monitor_outputs4,  // 监视输出4
    output reg [7:0] monitor_outputs5,  // 监视输出5
    output reg [7:0] monitor_outputs6,  // 监视输出6
    output reg [7:0] monitor_outputs7,  // 监视输出7
    output reg [7:0] monitor_outputs8,  // 监视输出8
    output reg [7:0] monitor_outputs9,  // 监视输出9
    output reg [7:0] monitor_outputs10, // 监视输出10
    output reg [7:0] monitor_outputs11, // 监视输出11
    output reg [7:0] monitor_outputs12, // 监视输出12
    output reg [7:0] monitor_outputs13, // 监视输出13
    output reg [7:0] monitor_outputs14, // 监视输出14
    output reg [7:0] monitor_outputs15  // 监视输出15
);
reg [7:0] memory [0:255];               // 16*16 = 256个8位机器码

initial begin
    // 这里可以预置一些机器码，作为初代版本
    memory[0] = 8'b00000001; // 示例机器码
    memory[1] = 8'b00000010; // 示例机器码
    memory[2] = 8'b00000011; // 示例机器码
    memory[3] = 8'b00000100; // 示例机器码
    // 可以继续填充其他机器码，直到memory[255]
end

always @(posedge clk) begin
    if (rst) begin
        opcode <= 32'b0;
    end else begin
        opcode <= {memory[(address+3)%256], memory[(address+2)%256], memory[(address+1)%256], memory[address]};
    end
end
always @(posedge clk) begin
    if (rst) begin
        monitor_outputs0 <= 8'b0;
        monitor_outputs1 <= 8'b0;
        monitor_outputs2 <= 8'b0;
        monitor_outputs3 <= 8'b0;
        monitor_outputs4 <= 8'b0;
        monitor_outputs5 <= 8'b0;
        monitor_outputs6 <= 8'b0;
        monitor_outputs7 <= 8'b0;
        monitor_outputs8 <= 8'b0;
        monitor_outputs9 <= 8'b0;
        monitor_outputs10 <= 8'b0;
        monitor_outputs11 <= 8'b0;
        monitor_outputs12 <= 8'b0;
        monitor_outputs13 <= 8'b0;
        monitor_outputs14 <= 8'b0;
        monitor_outputs15 <= 8'b0;
    end else begin
        monitor_outputs0 <= monitor_inputs0;
        monitor_outputs1 <= monitor_inputs1;
        monitor_outputs2 <= monitor_inputs2;
        monitor_outputs3 <= monitor_inputs3;
        monitor_outputs4 <= monitor_inputs4;
        monitor_outputs5 <= monitor_inputs5;
        monitor_outputs6 <= monitor_inputs6;
        monitor_outputs7 <= monitor_inputs7;
        monitor_outputs8 <= monitor_inputs8;
        monitor_outputs9 <= monitor_inputs9;
        monitor_outputs10 <= monitor_inputs10;
        monitor_outputs11 <= monitor_inputs11;
        monitor_outputs12 <= monitor_inputs12;
        monitor_outputs13 <= monitor_inputs13;
        monitor_outputs14 <= monitor_inputs14;
        monitor_outputs15 <= monitor_inputs15;
    end
end
endmodule
